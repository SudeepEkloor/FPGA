module three_bit_counter (
    input wire clk,
    input wire reset,  
    output reg [2:0] q
);

    always @(posedge clk) begin
        if (reset)
            q <= 3'b000;
        else
            q <= q + 1;
    end

endmodule
